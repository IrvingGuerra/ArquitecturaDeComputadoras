LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;
LIBRARY MACHXO2;
USE MACHXO2.ALL; 

ENTITY AND0 IS	PORT(
		AI00, BI00 : IN STD_LOGIC;
		AO00 : OUT STD_LOGIC
	);
END AND0;

ARCHITECTURE AND00 OF AND0 IS 
	BEGIN
		AO00<=AI00 AND BI00;
END ARCHITECTURE;
		