LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;
LIBRARY MACHXO2;
USE MACHXO2.ALL;
USE pakaguecom00.ALL;

ENTITY TOPADDER0 IS
	PORT(
		A0, B0 : in std_logic;
		S0, C0 : out std_logic
	);
END TOPADDER0;

ARCHITECTURE TOPADDER00 OF TOPADDER0 IS
BEGIN
	
	US000 : AND0 PORT MAP(
				AI00=>A0, 
				BI00=>B0,
				AO00=>C0
			);	
		
	US100 : XOR0 PORT MAP(
				AI00=>A0,
				BI00=>B0,
				AO00=>S0
			);
END TOPADDER00;